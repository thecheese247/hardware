-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 12.1 Build 177 11/07/2012 SJ Web Edition"
-- CREATED		"Thu Jan 17 19:39:01 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dlock IS 
	PORT
	(
		RESET :  IN  STD_LOGIC;
		CLOCK :  IN  STD_LOGIC;
		DATA :  IN  STD_LOGIC;
		LOCK :  OUT  STD_LOGIC;
		ALARM :  OUT  STD_LOGIC
	);
END dlock;

ARCHITECTURE bdf_type OF dlock IS 

SIGNAL	D0 :  STD_LOGIC;
SIGNAL	D1 :  STD_LOGIC;
SIGNAL	D2 :  STD_LOGIC;
SIGNAL	notDATA :  STD_LOGIC;
SIGNAL	notQ0 :  STD_LOGIC;
SIGNAL	notQ1 :  STD_LOGIC;
SIGNAL	notQ2 :  STD_LOGIC;
SIGNAL	notRESET :  STD_LOGIC;
SIGNAL	Q0 :  STD_LOGIC;
SIGNAL	Q1 :  STD_LOGIC;
SIGNAL	Q2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_12 <= '1';
SYNTHESIZED_WIRE_13 <= '1';
SYNTHESIZED_WIRE_14 <= '1';



D2 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_4 <= notDATA AND notQ1;


SYNTHESIZED_WIRE_3 <= DATA AND SYNTHESIZED_WIRE_7;


SYNTHESIZED_WIRE_7 <= Q0 OR Q2;


SYNTHESIZED_WIRE_6 <= Q2 AND Q0;


SYNTHESIZED_WIRE_5 <= notQ2 AND Q1 AND notQ0;


D0 <= SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_11 AND notQ2;


SYNTHESIZED_WIRE_8 <= DATA AND notQ1;


SYNTHESIZED_WIRE_2 <= Q1 AND Q0;


SYNTHESIZED_WIRE_9 <= Q2 AND Q0;


SYNTHESIZED_WIRE_11 <= DATA OR notQ0;


ALARM <= Q2 AND Q1 AND Q0;


PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_12)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_20 <= '0';
ELSIF (SYNTHESIZED_WIRE_12 = '0') THEN
	SYNTHESIZED_WIRE_20 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_20 <= D0;
END IF;
END PROCESS;



PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_13)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_22 <= '0';
ELSIF (SYNTHESIZED_WIRE_13 = '0') THEN
	SYNTHESIZED_WIRE_22 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_22 <= D2;
END IF;
END PROCESS;



notDATA <= NOT(DATA);



notQ0 <= NOT(SYNTHESIZED_WIRE_20);



PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_14)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_21 <= '0';
ELSIF (SYNTHESIZED_WIRE_14 = '0') THEN
	SYNTHESIZED_WIRE_21 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_21 <= D1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_15 AND DATA;


notRESET <= NOT(RESET);



Q0 <= SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_20;



notQ1 <= NOT(SYNTHESIZED_WIRE_21);



Q1 <= SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_21;


notQ2 <= NOT(SYNTHESIZED_WIRE_22);



Q2 <= SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_22;


LOCK <= NOT(Q2 AND Q1 AND notQ0);


SYNTHESIZED_WIRE_1 <= notQ1 AND SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_15 <= Q0 OR Q1;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_17 OR Q2;


SYNTHESIZED_WIRE_17 <= notDATA AND notQ0;


D1 <= SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19;


END bdf_type;