-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 12.1 Build 177 11/07/2012 SJ Web Edition"
-- CREATED		"Sun Jan 20 16:47:06 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dlock IS 
	PORT
	(
		RESET :  IN  STD_LOGIC;
		CLOCK :  IN  STD_LOGIC;
		DATA :  IN  STD_LOGIC;
		LOCK :  OUT  STD_LOGIC;
		ALARM :  OUT  STD_LOGIC
	);
END dlock;

ARCHITECTURE bdf_type OF dlock IS 

SIGNAL	D0 :  STD_LOGIC;
SIGNAL	D1 :  STD_LOGIC;
SIGNAL	D2 :  STD_LOGIC;
SIGNAL	notDATA :  STD_LOGIC;
SIGNAL	notQ0 :  STD_LOGIC;
SIGNAL	notQ1 :  STD_LOGIC;
SIGNAL	notQ2 :  STD_LOGIC;
SIGNAL	notRESET :  STD_LOGIC;
SIGNAL	Q0 :  STD_LOGIC;
SIGNAL	Q1 :  STD_LOGIC;
SIGNAL	Q2 :  STD_LOGIC;
SIGNAL	Q2norQ0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '1';
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_2 <= '1';



ALARM <= NOT(notQ2 OR notQ1 OR notQ0);


PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_0)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_19 <= '0';
ELSIF (SYNTHESIZED_WIRE_0 = '0') THEN
	SYNTHESIZED_WIRE_19 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_19 <= D0;
END IF;
END PROCESS;



PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_1)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_21 <= '0';
ELSIF (SYNTHESIZED_WIRE_1 = '0') THEN
	SYNTHESIZED_WIRE_21 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_21 <= D2;
END IF;
END PROCESS;



notDATA <= NOT(DATA);



notQ0 <= NOT(SYNTHESIZED_WIRE_19);



PROCESS(CLOCK,notRESET,SYNTHESIZED_WIRE_2)
BEGIN
IF (notRESET = '0') THEN
	SYNTHESIZED_WIRE_20 <= '0';
ELSIF (SYNTHESIZED_WIRE_2 = '0') THEN
	SYNTHESIZED_WIRE_20 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	SYNTHESIZED_WIRE_20 <= D1;
END IF;
END PROCESS;


notRESET <= NOT(RESET);



Q0 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_19;



notQ1 <= NOT(SYNTHESIZED_WIRE_20);



Q1 <= SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_20;


notQ2 <= NOT(SYNTHESIZED_WIRE_21);



Q2 <= SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_21;


D0 <= NOT(SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_5);


LOCK <= NOT(Q2 AND Q1 AND notQ0);


D2 <= NOT(SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_7 AND SYNTHESIZED_WIRE_8);


SYNTHESIZED_WIRE_4 <= NOT(notQ1 AND DATA);


SYNTHESIZED_WIRE_3 <= NOT(notQ2 AND SYNTHESIZED_WIRE_9);


SYNTHESIZED_WIRE_5 <= NOT(Q2norQ0);



SYNTHESIZED_WIRE_9 <= NOT(notDATA AND Q0);


D1 <= NOT(SYNTHESIZED_WIRE_10 AND SYNTHESIZED_WIRE_11);


SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13);


SYNTHESIZED_WIRE_10 <= NOT(SYNTHESIZED_WIRE_14 OR Q2norQ0);


SYNTHESIZED_WIRE_13 <= NOT(Q1 OR DATA);


SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_15 OR notDATA);


SYNTHESIZED_WIRE_15 <= NOT(Q0 OR Q2);


Q2norQ0 <= NOT(notQ0 OR notQ2);


SYNTHESIZED_WIRE_6 <= NOT(Q0 AND Q1);


SYNTHESIZED_WIRE_14 <= NOT(Q2 OR notQ1 OR Q0);


SYNTHESIZED_WIRE_7 <= NOT(DATA AND SYNTHESIZED_WIRE_16);


SYNTHESIZED_WIRE_8 <= NOT(SYNTHESIZED_WIRE_17 AND notQ1);


SYNTHESIZED_WIRE_16 <= NOT(notQ0 AND notQ1);


SYNTHESIZED_WIRE_17 <= NOT(SYNTHESIZED_WIRE_18 AND notQ2);


SYNTHESIZED_WIRE_18 <= NOT(notQ0 AND notDATA);


END bdf_type;